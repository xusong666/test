<<<<<<< HEAD
the first content is created by virtual machine 
the content is created by main laptop
=======
he first content is created by virtual machin
the second content is create by man bvir machine
the thirth content is created by loc bran vir mac
>>>>>>> 6ce03cc5ba2317294eefcb05b12927c863daa5c5
