the first content is created by virtual machine 

the content is created by loc bran vir mac
