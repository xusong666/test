the first content is created by virtual machine 
