he first content is created by virtual machin
the second content is create by man bvir machine
